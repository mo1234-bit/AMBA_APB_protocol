module test();
reg PCLK,PRESETn,transfer,READ_WRITE;
reg [8:0] apb_write_paddr;
reg [7:0]apb_write_data;
reg [8:0] apb_read_paddr;
wire PSLVERR;
wire [7:0] apb_read_data_out;
APB dut(PCLK,PRESETn,transfer,READ_WRITE,apb_write_paddr,apb_write_data,apb_read_paddr,PSLVERR,apb_read_data_out);
initial begin 
PCLK=0;
forever #1 PCLK=~PCLK;
end
initial begin 
PRESETn=0;
transfer=0;
READ_WRITE=0;
@(negedge PCLK);
PRESETn=1;
@(negedge PCLK);
transfer=1;
@(negedge PCLK);
@(negedge PCLK);
apb_write_paddr={1'b1,8'd60};
apb_write_data=8'b11011001;
@(negedge PCLK);
@(negedge PCLK);
apb_write_paddr={1'b1,8'd54};
apb_write_data=8'b10011101;
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
apb_write_paddr={1'b1,8'd43};
apb_write_data=8'b01011001;
@(negedge PCLK);
@(negedge PCLK);
apb_write_paddr={1'b1,8'd32};
apb_write_data=8'b10010001;
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
apb_write_paddr={1'b0,8'd12};
apb_write_data=8'b11111001;
@(negedge PCLK);
@(negedge PCLK);
apb_write_paddr={1'b0,8'd63};
apb_write_data=8'b10111011;
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
apb_write_paddr={1'b0,8'd34};
apb_write_data=8'b00111011;
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
apb_write_paddr={1'b0,8'd23};
apb_write_data=8'b10110011;
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
apb_write_paddr = 9'd526;
apb_write_data = 9'd9;
@(negedge PCLK);
@(negedge PCLK); 
apb_write_paddr = 9'd22; 
apb_write_data = 9'd23;
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
READ_WRITE=1;
PRESETn=0;
transfer=0;
@(negedge PCLK);
PRESETn=1;
@(negedge PCLK);
transfer=1;
apb_read_paddr={1'b1,8'd60};
@(negedge PCLK);
@(negedge PCLK);
apb_read_paddr={1'b1,8'd54};
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
apb_read_paddr={1'b1,8'd43};
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
apb_read_paddr={1'b1,8'd32};
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
apb_read_paddr={1'b0,8'd12};
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
apb_read_paddr={1'b0,8'd63};
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
apb_read_paddr={1'b0,8'd34};
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
apb_read_paddr={1'b0,8'd23};
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
apb_read_paddr={1'b0,8'b11011110};
@(negedge PCLK);
@(negedge PCLK);
@(negedge PCLK);
$stop;
end
endmodule
