module test();
reg PCLK,PRESETn,transfer,READ_WRITE;
reg [8:0] apb_write_paddr;
reg [7:0]apb_write_data;
reg [8:0] apb_read_paddr;
wire PSLVERR;
wire [7:0] apb_read_data_out;
APB dut(PCLK,PRESETn,transfer,READ_WRITE,apb_write_paddr,apb_write_data,apb_read_paddr,PSLVERR,apb_read_data_out);
initial begin 
PCLK=0;
forever #1 PCLK=~PCLK;
end
initial begin 
PRESETn=0;
transfer=0;
READ_WRITE=0;
@(negedge PCLK);
PRESETn=1;
@(negedge PCLK);
transfer=1;
repeat(2)@(negedge PCLK);
//@(negedge PCLK);
apb_write_paddr={1'b1,8'd60};
apb_write_data=8'b11011001;
repeat(2)@(negedge PCLK);
//@(negedge PCLK);
apb_write_paddr={1'b1,8'd54};
apb_write_data=8'b10011101;
repeat(5)@(negedge PCLK);
// @(negedge PCLK);
// @(negedge PCLK);
// @(negedge PCLK);
// @(negedge PCLK);
apb_write_paddr={1'b1,8'd43};
apb_write_data=8'b01011001;
repeat(2)@(negedge PCLK);
// @(negedge PCLK);
apb_write_paddr={1'b1,8'd32};
apb_write_data=8'b10010001;
repeat(3)@(negedge PCLK);
// @(negedge PCLK);
// @(negedge PCLK);
apb_write_paddr={1'b0,8'd12};
apb_write_data=8'b11111001;
repeat(2)@(negedge PCLK);
// @(negedge PCLK);
apb_write_paddr={1'b0,8'd63};
apb_write_data=8'b10111011;
repeat(3)@(negedge PCLK);
// @(negedge PCLK);
// @(negedge PCLK);
apb_write_paddr={1'b0,8'd34};
apb_write_data=8'b00111011;
repeat(4)@(negedge PCLK);
// @(negedge PCLK);
// @(negedge PCLK);
// @(negedge PCLK);
apb_write_paddr={1'b0,8'd23};
apb_write_data=8'b10110011;
repeat(6)@(negedge PCLK);
// @(negedge PCLK);
// @(negedge PCLK);
// @(negedge PCLK);
// @(negedge PCLK);
// @(negedge PCLK);
apb_write_paddr = 9'd526;
apb_write_data = 9'd9;
repeat(2)@(negedge PCLK);
// @(negedge PCLK); 
apb_write_paddr = 9'd22; 
apb_write_data = 9'd23;
repeat(4)@(negedge PCLK);
// @(negedge PCLK);
// @(negedge PCLK);
// @(negedge PCLK);
READ_WRITE=1;
PRESETn=0;
transfer=0;
@(negedge PCLK);
PRESETn=1;
@(negedge PCLK);
transfer=1;
apb_read_paddr={1'b1,8'd60};
repeat(2)@(negedge PCLK);
//@(negedge PCLK);
apb_read_paddr={1'b1,8'd54};
repeat(3)@(negedge PCLK);
//@(negedge PCLK);
//@(negedge PCLK);
apb_read_paddr={1'b1,8'd43};
repeat(3)@(negedge PCLK);
//@(negedge PCLK);
//@(negedge PCLK);
apb_read_paddr={1'b1,8'd32};
repeat(3)@(negedge PCLK);
//@(negedge PCLK);
//@(negedge PCLK);
apb_read_paddr={1'b0,8'd12};
repeat(3)@(negedge PCLK);
//@(negedge PCLK);
//@(negedge PCLK);
apb_read_paddr={1'b0,8'd63};
repeat(3)@(negedge PCLK);
//@(negedge PCLK);
//@(negedge PCLK);
apb_read_paddr={1'b0,8'd34};
repeat(3)@(negedge PCLK);
//@(negedge PCLK);
//@(negedge PCLK);
apb_read_paddr={1'b0,8'd23};
repeat(3)@(negedge PCLK);
//@(negedge PCLK);
//@(negedge PCLK);
apb_read_paddr={1'b0,8'b11011110};
repeat(3)@(negedge PCLK);
//@(negedge PCLK);
//@(negedge PCLK);
$stop;
end
endmodule
